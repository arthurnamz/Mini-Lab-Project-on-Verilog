`timescale 1ns/1ps

module memory_tb;



endmodule